/*
 * This module performs the shifting operations 
 */ 

module shift(input logic [6:0] sh,
				 input logic [31:0] RD2,
				 output logic [31:0] y);
	
	// AQUI DEBEN IR LAS OPERACIONES DE SHIFT
	
	always_comb
	
	
endmodule
